`timescale 1ns / 1ps
module lab4_b_tb;

  reg [3:0] a, b, c, d;
  reg [2:0] x, y, z;
  wire A, B, C, D, E, F, G, s1, s2, s3, s4, s5, s6, s7, s8, DP;

  lab4_b dut (
    .a(a),
    .b(b),
    .c(c),
    .d(d),
    .x(x),
    .y(y),
    .z(z),
    .A(A),
    .B(B),
    .C(C),
    .D(D),
    .E(E),
    .F(F),
    .G(G),
    .s1(s1),
    .s2(s2),
    .s3(s3),
    .s4(s4),
    .s5(s5),
    .s6(s6),
    .s7(s7),
    .s8(s8),
    .DP(DP)
  );

  initial begin
    $dumpfile("dump.vcd");
    $dumpvars(0, lab4_b_tb, A, B, C, D, E, F, G, DP, s1, s2, s3, s4, s5, s6, s7, s8);
    a = 4'b0000; b = 4'b0000; c = 4'b0000; d = 4'b0000;
    x = 3'b000; y = 3'b000; z = 3'b000;
    #10;

    // Case 0001
    a = 4'b0000; b = 4'b0000; c = 4'b0000; d = 4'b0001;
    x = 3'b000; y = 3'b000; z = 3'b001;
    #10;

    // Case 0010
    a = 4'b0000; b = 4'b0000; c = 4'b0001; d = 4'b0000;
    x = 3'b000; y = 3'b001; z = 3'b000;
    #10;

    // Case 0011
    a = 4'b0000; b = 4'b0000; c = 4'b0001; d = 4'b0001;
    x = 3'b000; y = 3'b001; z = 3'b001;
    #10;

    // Case 0100
    a = 4'b0000; b = 4'b0001; c = 4'b0000; d = 4'b0000;
    x = 3'b000; y = 3'b010; z = 3'b000;
    #10;

    // Case 0101
    a = 4'b0000; b = 4'b0001; c = 4'b0000; d = 4'b0001;
    x = 3'b000; y = 3'b010; z = 3'b001;
    #10;

    // Case 0110
    a = 4'b0000; b = 4'b0001; c = 4'b0001; d = 4'b0000;
    x = 3'b000; y = 3'b011; z = 3'b000;
    #10;

    // Case 0111
    a = 4'b0000; b = 4'b0001; c = 4'b0001; d = 4'b0001;
    x = 3'b000; y = 3'b011; z = 3'b001;
    #10;

    // Case 1000
    a = 4'b0001; b = 4'b0000; c = 4'b0000; d = 4'b0000;
    x = 3'b001; y = 3'b000; z = 3'b000;
    #10;

    // Case 1001
    a = 4'b0001; b = 4'b0000; c = 4'b0000; d = 4'b0001;
    x = 3'b001; y = 3'b000; z = 3'b001;
    #10;

    // Case 1010
    a = 4'b0001; b = 4'b0000; c = 4'b0001; d = 4'b0000;
    x = 3'b001; y = 3'b001; z = 3'b000;
    #10;

    // Case 1011
    a = 4'b0001; b = 4'b0000; c = 4'b0001; d = 4'b0001;
    x = 3'b001; y = 3'b001; z = 3'b001;
    #10;

    // Case 1100
    a = 4'b0001; b = 4'b0001; c = 4'b0000; d = 4'b0000;
    x = 3'b001; y = 3'b010; z = 3'b000;
    #10;

    // Case 1101
    a = 4'b0001; b = 4'b0001; c = 4'b0000; d = 4'b0001;
    x = 3'b001; y = 3'b010; z = 3'b001;
    #10;

    // Case 1110
    a = 4'b0001; b = 4'b0001; c = 4'b0001; d = 4'b0000;
    x = 3'b001; y = 3'b011; z = 3'b000;
    #10;

    // Case 1111
    a = 4'b0001; b = 4'b0001; c = 4'b0001; d = 4'b0001;
    x = 3'b001; y = 3'b011; z = 3'b001;
    #10;

    // Test Cases for xyz
    // Case 000
    a = 4'b0000; b = 4'b0000; c = 4'b0000; d = 4'b0000;
    x = 3'b000; y = 3'b000; z = 3'b000;
    #10;

    // Case 001
    a = 4'b0000; b = 4'b0000; c = 4'b0000; d = 4'b0000;
    x = 3'b000; y = 3'b000; z = 3'b001;
    #10;

    // Case 010
    a = 4'b0000; b = 4'b0000; c = 4'b0000; d = 4'b0000;
    x = 3'b000; y = 3'b001; z = 3'b000;
    #10;

    // Case 011
    a = 4'b0000; b = 4'b0000; c = 4'b0000; d = 4'b0000;
    x = 3'b000; y = 3'b001; z = 3'b001;
    #10;

    // Case 100
    a = 4'b0000; b = 4'b0000; c = 4'b0000; d = 4'b0000;
    x = 3'b001; y = 3'b000; z = 3'b000;
    #10;

    // Case 101
    a = 4'b0000; b = 4'b0000; c = 4'b0000; d = 4'b0000;
    x = 3'b001; y = 3'b000; z = 3'b001;
    #10;

    // Case 110
    a = 4'b0000; b = 4'b0000; c = 4'b0000; d = 4'b0000;
    x = 3'b001; y = 3'b001; z = 3'b000;
    #10;

    // Case 111
    a = 4'b0000; b = 4'b0000; c = 4'b0000; d = 4'b0000;
    x = 3'b001; y = 3'b001; z = 3'b001;
    #10;

    // End simulation
    $finish;
  end

endmodule
